module vga_clock(clk, clock_out);

	// Señal de reloj de entrada proveniente del FPGA
	input clk;
	
	// Señal de reloj de salida después de dividir la frecuencia
	output reg clock_out;

	// Registro de 28 bits que cuenta el número de ciclos de reloj de entrada
	reg[27:0] counter = 28'd0;
	
	// Valor por el cual se dividirá la frecuencia de la señal de entrada
	parameter DIVISOR = 28'd5000000;
	
	// The frequency of the output clk_out
	//  = The frequency of the input clk_in divided by DIVISOR
	// For example: Fclk_in = 50Mhz, if you want to get 1Hz signal to blink LEDs
	// You will modify the DIVISOR parameter value to 28'd50.000.000
	// Then the frequency of the output clk_out = 50Mhz/50.000.000 = 1Hz
	
	always @(posedge clk) begin
		counter <= counter + 28'd1;
			if (counter >= (DIVISOR-1))
				counter <= 28'd0;
		clock_out <= (counter < DIVISOR/2) ? 1'b1 : 1'b0;
	end
	
endmodule