module regressiveCounter(input wire [N-1:0] binary_input,
								 output wire [N-1:0] binary_output);

	assign binary_output = binary_input - 1;

endmodule